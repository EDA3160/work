.SUBCKT AN2D2 A1 A2 Z VDD VSS
MM9 net14 A2 VSS VSS nch_mac l=30.0n w=0.14u
MM8 net26 A1 net14 VSS nch_mac l=30.0n w=0.14u
MM5 Z net26 VSS VSS nch_mac l=30.0n w=0.14u
MM5_2 Z net26 VSS VSS nch_mac l=30.0n w=0.14u
MM6 net26 A1 VDD VDD pch_mac l=30.0n w=170.0n
MM7 net26 A2 VDD VDD pch_mac l=30.0n w=0.17u
MM4 Z net26 VDD VDD pch_mac l=30.0n w=0.17u
MM4_2 Z net26 VDD VDD pch_mac l=30.0n w=0.17u
.ENDS